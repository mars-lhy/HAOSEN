------------------------------------------------------------------------
-- effects_layer.vhd
------------------------------------------------------------------------
-- Author : Ulrich Zolt�n
--          Copyright 2006 Digilent, Inc.
------------------------------------------------------------------------
-- Software version : Xilinx ISE 7.1.04i
--                    WebPack
-- Device	        : 3s200ft256-4
------------------------------------------------------------------------
-- This file describes logic to make the negative and grayscale effects
-- on the incoming pixels in real time, effect being selected by input
-- from the keyboard_controller. Both negative and grayscale can be
-- applied at the same time. Effects are applied only while inside the
-- image boundaries, the rest of the pixels pass unaltered.
------------------------------------------------------------------------
--  Behavioral description
------------------------------------------------------------------------
-- The 3 color channel, each 4 bits width, generated by the
-- image_controller are inputs to this module. The image_controller also
-- generates the input inside_image which is active when current pixel
-- is contained in the image and is not part of the background.
-- The keyboard send the last generated ascii character, together with
-- event_type signal and new_key, active for one clock period when a new
-- key event is generated. event_type is low when a key was pressed on
-- the keyboard, or it was held down. This is called a MAKE event.
-- event_type is high when a key was released, BREAK event.
-- To activate negative effect, the N key must be pressed (MAKE event on
--  N key). Another MAKE event on N key will disable the negative effect
-- Similar to the negative, grayscale effect can be toggled by pressing
-- G key.
-- Making the negative of the image is easily done by xor-ing the pixel
-- data with 1 (4 bits of 1), which is equivalent to inverting the pixel
-- For the grayscale effect, a gray intensity is computed by multipling
-- each color channel with a weight(dependant on the wave length of the
-- corresponding channel) and the results are added to obtain the gray
-- intensity. This intensity is attributed to each color channel.
-- The weights are: 0.30 for red
--                  0.58 for green; human eye is more sensitive to green
--                  0.12 for blue
-- For making this multiplications, the values of the channels received
-- from the image_controller is multiplied by an integer (using the
-- multipliers on the spartan3 fpga), added and the result is shifted
-- 9 bits to the right, which is equivalent to (integer) division by 512
-- The integers used for multipling are:
-- 154 for red  : 154/512 = 0.30078125
-- 298 for green: 298/512 = 0.58203125
--  60 for blue :  60/512 = 0.11718750
-- 154 + 298 + 60 = 512, otherwise image luminosity would be altered
------------------------------------------------------------------------
--  Port definitions
------------------------------------------------------------------------
-- clk         - global clock input of 100MHz
-- red_in      - red channel data of the pixel from image_controller
-- green_in    - green channel data of the pixel from image_controller
-- blue_in     - blue channel data of the pixel from image_controller
-- inside_image- input pin from image_controller, high when pixel is
--             - part of the image, else pixel is from background
-- ascii_in    - input, 7 bits, from keyboard_controller, indicates
--             - ascii code of last pressed key.
-- event_type  - input, from keyboard controller, low when last event
--             - was a MAKE event, high when it was a BREAK event
-- new_key     - input, from keyboard_controller, indicates a new event
--             - occurred and ascii code and event type is valid on
--             - ascii_in and event_type respectively
-- red_out     - output, 4 bits, red color channel of the altered pixel
--             - if any effect were applied to it, else it is the same
--             - as red_in
-- green_out   - output, 4 bits, green color channel of the altered
--             - pixel if any effect were applied to it, else it is the
--             - same as green_in
-- blue_out    - output, 4 bits, blue color channel of the altered pixel
--             - if any effect were applied to it, else it is the same
--             - as blue_in
------------------------------------------------------------------------
-- Revision History:
-- 09/18/2006(UlrichZ): created
------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- simulation library
library UNISIM;
use UNISIM.VComponents.all;

-- the effects_layer entity declaration
-- read above for behavioral description and port definitions.
entity effects_layer is
port(
   clk         : in std_logic;

   red_in      : in std_logic_vector(3 downto 0);
   green_in    : in std_logic_vector(3 downto 0);
   blue_in     : in std_logic_vector(3 downto 0);
   inside_image: in std_logic;

   ascii_in    : in std_logic_vector(6 downto 0);
   event_type  : in std_logic;
   new_key     : in std_logic;

   red_out     : out std_logic_vector(3 downto 0);
   green_out   : out std_logic_vector(3 downto 0);
   blue_out    : out std_logic_vector(3 downto 0)
);
end effects_layer;

architecture Behavioral of effects_layer is

------------------------------------------------------------------------
-- SIGNALS
------------------------------------------------------------------------

-- active when negative effect should be applied
signal negative_on  : std_logic := '0';
-- active when grayscale effect should be applied
signal grayscale_on : std_logic := '0';

------------------------------------------------------------------------
-- CONSTANTS
------------------------------------------------------------------------

constant LETTER_N : std_logic_vector(6 downto 0) := "1101110"; -- 0x6E
constant LETTER_G : std_logic_vector(6 downto 0) := "1100111"; -- 0x67
constant MAKE_EVENT : std_logic := '0';

-- the integer weights represented on 9 bits
constant N_154 : std_logic_vector(8 downto 0) := "010011010";  -- 154
constant N_298 : std_logic_vector(8 downto 0) := "100101010";  -- 298
constant N_060 : std_logic_vector(8 downto 0) := "000111100";  --  60

begin

   -- this process applies the effects on the incoming pixels
   -- uses variable to store intermediary results
   -- first applies the grayscale effect if needed, then
   -- the negative (also if needed)
   process(clk)
   -- hold the result of the multiplication of the red channel value
   -- with the corresponding integer weight
   variable product_red  : std_logic_vector(12 downto 0);
   -- hold the result of the multiplication of the green channel value
   -- with the corresponding integer weight   
   variable product_green: std_logic_vector(12 downto 0);
   -- hold the result of the multiplication of the blue channel value
   -- with the corresponding integer weight
   variable product_blue : std_logic_vector(12 downto 0);
   -- value of the gray intensity obtained by adding the above products
   -- and shifting the result 9 bits to the right (division by 512).
   variable gray : std_logic_vector(12 downto 0);
   -- intermediary values for the output color channels
   variable temp_red  : std_logic_vector(3 downto 0);
   variable temp_green: std_logic_vector(3 downto 0);
   variable temp_blue : std_logic_vector(3 downto 0);
   begin
      if(rising_edge(clk)) then
         -- if pixel is part of the image
         if(inside_image = '1') then
            -- assign original values
            temp_red := red_in;
            temp_green := green_in;
            temp_blue := blue_in;
            -- if the grayscale should be applied
            if(grayscale_on = '1') then
               -- make the multiplications
               product_red   := red_in * N_154;
               product_green := green_in * N_298;
               product_blue  := blue_in * N_060;
               -- add the products
               gray := product_red + product_green + product_blue;
               -- make the division by 512 and assing gray intensity
               -- to color channels
               temp_red   := gray(12 downto 9);
               temp_green := gray(12 downto 9);
               temp_blue  := gray(12 downto 9);
            end if;
            -- if the negative should be applied
            -- Notice else keyword is nit used, because both
            -- effect could be applied simultaneously
            -- This is the reason for using variables instead of signals
            if(negative_on = '1') then
               -- xor the channel value with 1 to invert the value
               temp_red   := temp_red xor "1111";
               temp_green := temp_green xor "1111";
               temp_blue  := temp_blue xor "1111";
            end if;
            -- assign intermediary values to outputs
            red_out <= temp_red;
            green_out <= temp_green;
            blue_out <= temp_blue;
         else
            -- no effect should be applied to the background
            red_out <= red_in;
            green_out <= green_in;
            blue_out <= blue_in;
         end if;
      end if;
   end process;

   -- checks for new key event, and if MAKE event and letter N pressed
   -- then set negative_on high. Similarly for grayscale is G is pressed
   process(clk)
   begin
      if(rising_edge(clk)) then
         if(new_key = '1' and event_type = MAKE_EVENT) then
            if(ascii_in = LETTER_N) then
               negative_on <= not negative_on;
            elsif(ascii_in = LETTER_G) then
               grayscale_on <= not grayscale_on;
            end if;
         end if;
      end if;
   end process;

end Behavioral;
