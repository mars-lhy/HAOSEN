library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity DigitalSynth is
	port (
		clk			: in STD_LOGIC; -- Master clock (50 MHz)
		rst			: in STD_LOGIC; -- Reset button (synchronous reset)
		kd				: in STD_LOGIC; -- PS/2 keyboard data signal
		kc				: in STD_LOGIC; -- PS/2 keyboard clock signal
		sclk			: out STD_LOGIC; -- Serial clock of the DAC (Digital-to-Analog Converter)
		sync			: out STD_LOGIC; -- Synchronize signal
		sdata			: out STD_LOGIC; -- Serial data
		eppDataBus	: inout STD_LOGIC_VECTOR(7 downto 0); -- EPP protocol data bus
		eppAstb		: in STD_LOGIC; -- EPP protocol address strobe
		eppDstb		: in STD_LOGIC; -- EPP protocol data strobe
		eppWrite		: in STD_LOGIC; -- EPP protocol write signal
		eppWait		: out STD_LOGIC -- EPP protocol wait signal
	);
end DigitalSynth;

architecture Behavioral of DigitalSynth is

	-- This component handles the keyboard operation, including the polyphony arbitration.
	component KeyboardUnit is
		port (
			clk		: in STD_LOGIC;
			rst		: in STD_LOGIC;
			kc			: in STD_LOGIC;
			kd			: in STD_LOGIC;
			kbNote0	: out STD_LOGIC_VECTOR(4 downto 0);
			kbNote1	: out STD_LOGIC_VECTOR(4 downto 0);
			kbNote2	: out STD_LOGIC_VECTOR(4 downto 0);
			kbNote3	: out STD_LOGIC_VECTOR(4 downto 0);
			kbStatus	: out STD_LOGIC_VECTOR(3 downto 0)
		);
	end component;

	-- This component handles the USB communication (the EPP protocol).
	component UsbUnit is
		port (
			clk				: in STD_LOGIC;
			eppAstb			: in STD_LOGIC;
			eppDstb			: in STD_LOGIC;
			eppWrite			: in STD_LOGIC;
			eppWait			: out STD_LOGIC;
			eppDataBus		: inout STD_LOGIC_VECTOR(7 downto 0);
			usbNote0			: out STD_LOGIC_VECTOR(4 downto 0);
			usbNote1			: out STD_LOGIC_VECTOR(4 downto 0);
			usbNote2			: out STD_LOGIC_VECTOR(4 downto 0);
			usbNote3			: out STD_LOGIC_VECTOR(4 downto 0);
			usbStatus		: out STD_LOGIC_VECTOR(3 downto 0);
			midiDirection	: in STD_LOGIC;
			midiNote0		: in STD_LOGIC_VECTOR(4 downto 0);
			midiNote1		: in STD_LOGIC_VECTOR(4 downto 0);
			midiNote2		: in STD_LOGIC_VECTOR(4 downto 0);
			midiNote3		: in STD_LOGIC_VECTOR(4 downto 0);
			midiStatus		: in STD_LOGIC_VECTOR(3 downto 0);
			control			: out STD_LOGIC_VECTOR(7 downto 0);
			parameter0		: out STD_LOGIC_VECTOR(7 downto 0);
			parameter1		: out STD_LOGIC_VECTOR(7 downto 0);
			parameter2		: out STD_LOGIC_VECTOR(7 downto 0);
			parameter3		: out STD_LOGIC_VECTOR(7 downto 0)
		);
	end component;

	-- This component select between the notes and status generated by the keyboard
	-- and those received via USB. The chosen notes and status drives the oscillators.
	component NoteSelector is
		port (
			selector											: in STD_LOGIC;
			kbNote0, kbNote1, kbNote2, kbNote3		: in STD_LOGIC_VECTOR(4 downto 0);
			usbNote0, usbNote1, usbNote2, usbNote3	: in STD_LOGIC_VECTOR(4 downto 0);
			note0, note1, note2, note3					: out STD_LOGIC_VECTOR(4 downto 0);
			kbStatus											: in STD_LOGIC_VECTOR(3 downto 0);
			usbStatus										: in STD_LOGIC_VECTOR(3 downto 0);
			status											: out STD_LOGIC_VECTOR(3 downto 0)
		);
	end component;

	-- This component represents the 4 oscillators (corresponding to the 4-note polyphony).
	component OscillatorsUnit is
		port (
			clk					: in STD_LOGIC;
			rst					: in STD_LOGIC;
			waveType				: in STD_LOGIC;
			oscillatorStatus	: in STD_LOGIC_VECTOR(3 downto 0);
			noteAddress0		: in STD_LOGIC_VECTOR(4 downto 0);
			noteAddress1		: in STD_LOGIC_VECTOR(4 downto 0);
			noteAddress2		: in STD_LOGIC_VECTOR(4 downto 0);
			noteAddress3		: in STD_LOGIC_VECTOR(4 downto 0);
			outputWave			: out STD_LOGIC_VECTOR(7 downto 0)
		);
	end component;

	-- This component applies audio effects to the waves generated by the oscillators.
	component EffectsUnit is
		port (
			clk				: in STD_LOGIC;
			effectSelect	: in STD_LOGIC_VECTOR(1 downto 0);
			parameter		: in STD_LOGIC_VECTOR(7 downto 0);
			feedbackAmount	: in STD_LOGIC_VECTOR(7 downto 0);
			wetAmount		: in STD_LOGIC_VECTOR(7 downto 0);
			dryAmount		: in STD_LOGIC_VECTOR(7 downto 0);
			originalData	: in STD_LOGIC_VECTOR(7 downto 0);
			processedData	: out STD_LOGIC_VECTOR(7 downto 0)
		);
	end component;

	-- This component sends serialized data to the digital-to-analog converter.
	component SpiUnit is
		port (
			clk		: in STD_LOGIC;
			data		: in STD_LOGIC_VECTOR(7 downto 0);
			control	: in STD_LOGIC_VECTOR(7 downto 0);
			sclk		: out STD_LOGIC;
			sync		: out STD_LOGIC;
			sdata		: out STD_LOGIC
		);
	end component;

	signal kbNote0, kbNote1, kbNote2, kbNote3			: STD_LOGIC_VECTOR(4 downto 0);
	signal usbNote0, usbNote1, usbNote2, usbNote3	: STD_LOGIC_VECTOR(4 downto 0);
	signal note0, note1, note2, note3					: STD_LOGIC_VECTOR(4 downto 0);
	signal kbStatus, usbStatus, status					: STD_LOGIC_VECTOR(3 downto 0);

	signal spiData, outputWave								: STD_LOGIC_VECTOR(7 downto 0);
	signal param0, param1, param2, param3, control	: STD_LOGIC_VECTOR(7 downto 0);

begin

	KeyboardUnit_Map: KeyboardUnit port map (
		clk => clk,
		rst => rst,
		kc => kc,
		kd => kd,
		kbNote0 => kbNote0,
		kbNote1 => kbNote1,
		kbNote2 => kbNote2,
		kbNote3 => kbNote3,
		kbStatus => kbStatus
	);

	UsbUnit_Map: UsbUnit port map (
		clk => clk,
		eppAstb => eppAstb,
		eppDstb => eppDstb,
		eppWrite => eppWrite,
		eppWait => eppWait,
		eppDataBus => eppDataBus,
		usbNote0 => usbNote0,
		usbNote1 => usbNote1,
		usbNote2 => usbNote2,
		usbNote3 => usbNote3,
		usbStatus => usbStatus,
		midiDirection => control(0),
		midiNote0 => kbNote0,
		midiNote1 => kbNote1,
		midiNote2 => kbNote2,
		midiNote3 => kbNote3,
		midiStatus => kbStatus,
		control => control,
		parameter0 => param0,
		parameter1 => param1,
		parameter2 => param2,
		parameter3 => param3
	);

	NoteSelector_Map: NoteSelector port map (
		selector => control(0),
		kbNote0 => kbNote0,
		kbNote1 => kbNote1,
		kbNote2 => kbNote2,
		kbNote3 => kbNote3,
		usbNote0 => usbNote0,
		usbNote1 => usbNote1,
		usbNote2 => usbNote2,
		usbNote3 => usbNote3,
		note0 => note0,
		note1 => note1,
		note2 => note2,
		note3 => note3,
		kbStatus => kbStatus,
		usbStatus => usbStatus,
		status => status
	);

	OscillatorsUnit_Map: OscillatorsUnit port map (
		clk => clk,
		rst => rst,
		waveType => control(7),
		oscillatorStatus => status,
		noteAddress0 => note0,
		noteAddress1 => note1,
		noteAddress2 => note2,
		noteAddress3 => note3,
		outputWave => outputWave
	);

	EffectsUnit_Map: EffectsUnit port map (
		clk => clk,
		effectSelect => control(2 downto 1),
		parameter => param0,
		feedbackAmount => param1,
		wetAmount => param2,
		dryAmount => param3,
		originalData => outputWave,
		processedData => spiData
	);

	SpiUnit_Map: SpiUnit port map (
		clk => clk,
		data => spiData,
		control => x"10",
		sclk => sclk,
		sync => sync,
		sdata => sdata
	);

end Behavioral;