------------------------------------------------------------------------
--	NoteSelector.vhd
------------------------------------------------------------------------
--	Author:	Lucian Chetan
------------------------------------------------------------------------
--	Software version: Xilinx WebPack ISE 8.1i
------------------------------------------------------------------------
--	The module selects between the notes and status generated by the keyboard unit
--	and the notes and status received by the USB unit. The signal that decides
--	the source of the notes and status comes from the USB unit, being controlled
--	by the software application. The keyboard is active only when the user records
--	a MIDI file or simply plays. When the user plays a MIDI file, the keyboard
--	is inactive, and the notes sent by the software application are rendered by
--	the oscillators.
------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity NoteSelector is
	port (
		selector											: in STD_LOGIC; -- '0' => keyboard notes, '1' => USB notes
		kbNote0, kbNote1, kbNote2, kbNote3		: in STD_LOGIC_VECTOR(4 downto 0); -- Data from the keyboard
		usbNote0, usbNote1, usbNote2, usbNote3	: in STD_LOGIC_VECTOR(4 downto 0); -- Data from the USB module
		note0, note1, note2, note3					: out STD_LOGIC_VECTOR(4 downto 0); -- Data to the oscillators
		kbStatus											: in STD_LOGIC_VECTOR(3 downto 0); -- Status from the keyboard
		usbStatus										: in STD_LOGIC_VECTOR(3 downto 0); -- Status from the USB module
		status											: out STD_LOGIC_VECTOR(3 downto 0) -- Status to the oscillators
	);
end NoteSelector;

architecture Behavioral of NoteSelector is

begin

	-- If "selector" = '0', then the source of the notes and status for the oscillators is the keyboard unit.
	-- If "selector" = '1', then the source of the notes and status for the oscillators is the USB unit.
	note0 <= kbNote0 when (selector = '0') else usbNote0;
	note1 <= kbNote1 when (selector = '0') else usbNote1;
	note2 <= kbNote2 when (selector = '0') else usbNote2;
	note3 <= kbNote3 when (selector = '0') else usbNote3;
	status <= kbStatus when (selector = '0') else usbStatus;
	
end Behavioral;