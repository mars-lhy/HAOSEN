------------------------------------------------------------------------
--	OscillatorGroup.vhd
------------------------------------------------------------------------
--	Author:	Lucian Chetan
------------------------------------------------------------------------
--	Software version: Xilinx WebPack ISE 8.1i
------------------------------------------------------------------------
--	This module groups the modules that:
--		-	generate a wave according to the note periods ("Oscillator"),
--		-	resample the data at 48 kHz ("Sampler").
------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity OscillatorGroup is
	port (
		clk					: in STD_LOGIC; -- Master clock (50 MHz)
		rst					: in STD_LOGIC; -- Reset button (synchronous reset)
		waveType				: in STD_LOGIC; -- The type of wave generated by the oscillators: '0' = sawtooth, '1'  = square
		oscillatorStatus	: in STD_LOGIC_VECTOR(3 downto 0); -- The status of the oscillators
		notePeriod0			: in STD_LOGIC_VECTOR(10 downto 0); -- The period of the first note
		notePeriod1			: in STD_LOGIC_VECTOR(10 downto 0); -- The period of the second note
		notePeriod2			: in STD_LOGIC_VECTOR(10 downto 0); -- The period of the third note
		notePeriod3			: in STD_LOGIC_VECTOR(10 downto 0); -- The period of the fourth note
		outputWave			: out STD_LOGIC_VECTOR(7 downto 0) -- The sum of all four waves
	);
end OscillatorGroup;

architecture Behavioral of OscillatorGroup is

	-- This component represents the oscillator whose waveform is enveloped using the ADSR amplitude modulation model.
	component Oscillator is
		port (
			clk					: in STD_LOGIC;
			rst					: in STD_LOGIC;
			waveType				: in STD_LOGIC;
			oscillatorStatus	: in STD_LOGIC;
			notePeriod			: in STD_LOGIC_VECTOR(10 downto 0);
			outputWave			: out STD_LOGIC_VECTOR(15 downto 0)
		);
	end component;
	
	-- This component represents the adder that adds the 4 waves generated by the 4 oscillators.
	component Adder is
		port (
			a			: in STD_LOGIC_VECTOR(15 downto 0);
			b			: in STD_LOGIC_VECTOR(15 downto 0);
			c			: in STD_LOGIC_VECTOR(15 downto 0);
			d			: in STD_LOGIC_VECTOR(15 downto 0);
			output	: out STD_LOGIC_VECTOR(7 downto 0)
		);
	end component;
	
	signal w0, w1, w2, w3: STD_LOGIC_VECTOR(15 downto 0);

begin

	Oscillator0_Map: Oscillator port map (
		clk => clk,
		rst => rst,
		waveType => waveType,
		oscillatorStatus => oscillatorStatus(0),
		notePeriod => notePeriod0,
		outputWave => w0
	);
	
	Oscillator1_Map: Oscillator port map (
		clk => clk,
		rst => rst,
		waveType => waveType,
		oscillatorStatus => oscillatorStatus(1),
		notePeriod => notePeriod1,
		outputWave => w1
	);
	
	Oscillator2_Map: Oscillator port map (
		clk => clk,
		rst => rst,
		waveType => waveType,
		oscillatorStatus => oscillatorStatus(2),
		notePeriod => notePeriod2,
		outputWave => w2
	);
	
	Oscillator3_Map: Oscillator port map (
		clk => clk,
		rst => rst,
		waveType => waveType,
		oscillatorStatus => oscillatorStatus(3),
		notePeriod => notePeriod3,
		outputWave => w3
	);
	
	Adder_Map: Adder port map (
		a => w0,
		b => w1,
		c => w2,
		d => w3,
		output => outputWave
	);

end Behavioral;