--------------------------------------------------------------------------------
-- Company: 
-- Author: Fazakas Szabolcs
--
-- Create Date:    00:02:49 10/05/06
-- Design Name:    
-- Module Name:    video - Behavioral
-- Project Name:   
-- Target Device:  
-- Tool versions:  
-- Description:
--
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
Library UNISIM;
use UNISIM.vcomponents.all;
---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
------------------------------------------------------------------------
-- This component has 4 BlockRams which contains the images for the 
-- video.
--
------------------------------------------------------------------------
--  Port definitions
------------------------------------------------------------------------
-- mclk             Input      Main clock input 
-- frame(15:0)      Input      Address
-- laser            Output     Data output
--
------------------------------------------------------------------------
entity video is
 Port(    mclk    : in std_logic;
          frame   : in std_logic_vector(15 downto 0);

        laser           :out std_logic
        );
end video;

architecture Behavioral of video is
------------------------------------------------------------------------
-- Component Declarations
------------------------------------------------------------------------

------------------------------------------------------------------------
-- Signal Declarations
------------------------------------------------------------------------

 signal addres1,addres2,addres3,addres4  : std_logic_vector(13 downto 0);
 signal pixel1,pixel2,pixel3,pixel4: std_logic_vector(0 downto 0);
 
------------------------------------------------------------------------
-- Module Implementation - 
------------------------------------------------------------------------

begin

    addres1<=frame(13 downto 0);
    addres2<=frame(13 downto 0);
    addres3<=frame(13 downto 0);
    addres4<=frame(13 downto 0);

    laser<=pixel1(0) when frame(15 downto 14)="00" else
           pixel2(0) when frame(15 downto 14)="01" else 
           pixel3(0) when frame(15 downto 14)="10" else
           pixel4(0) when frame(15 downto 14)="11" else
           '0';
  
  
  RAMB16_S1_inst1 : RAMB16_S1
   generic map (
      INIT => "0", --  Value of output RAM registers at startup
      SRVAL => "0", --  Ouput value upon SSR assertion
      WRITE_MODE => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_01 => X"8000000080000000800000008000000080000000800000008000000080000000",
INIT_02 => X"E0000000E0000000E0000000E0000000E0000000E0000000E0000000E0000000",
INIT_03 => X"F8000000F8000000F8000000F8000000F8000000F8000000F8000000F8000000",
INIT_04 => X"FE000000FE000000FE000000FE000000FE000000FE000000FE000000FE000000",
INIT_05 => X"FF800000FF800000FF800000FF800000FF800000FF800000FF800000FF800000",
INIT_06 => X"FFE00000FFE00000FFE00000FFE00000FFE00000FFE00000FFE00000FFE00000",
INIT_07 => X"FFF80000FFF80000FFF80000FFF80000FFF80000FFF80000FFF80000FFF80000",
INIT_08 => X"FFFE0000FFFE0000FFFE0000FFFE0000FFFE0000FFFE0000FFFE0000FFFE0000",
INIT_09 => X"FFFF8000FFFF8000FFFF8000FFFF8000FFFF8000FFFF8000FFFF8000FFFF8000",
INIT_0a => X"FFFFE000FFFFE000FFFFE000FFFFE000FFFFE000FFFFE000FFFFE000FFFFE000",
INIT_0b => X"FFFFF800FFFFF800FFFFF800FFFFF800FFFFF800FFFFF800FFFFF800FFFFF800",
INIT_0c => X"FFFFFE00FFFFFE00FFFFFE00FFFFFE00FFFFFE00FFFFFE00FFFFFE00FFFFFE00",
INIT_0d => X"FFFFFF80FFFFFF80FFFFFF80FFFFFF80FFFFFF80FFFFFF80FFFFFF80FFFFFF80",
INIT_0e => X"FFFFFFE0FFFFFFE0FFFFFFE0FFFFFFE0FFFFFFE0FFFFFFE0FFFFFFE0FFFFFFE0",
INIT_0f => X"FFFFFFF8FFFFFFF8FFFFFFF8FFFFFFF8FFFFFFF8FFFFFFF8FFFFFFF8FFFFFFF8",
INIT_10 => X"FFFFFFFEFFFFFFFEFFFFFFFEFFFFFFFEFFFFFFFEFFFFFFFEFFFFFFFEFFFFFFFE",
INIT_11 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_12 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_13 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_14 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_15 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_16 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
INIT_17 => X"1FFFFFFF1FFFFFFF1FFFFFFF1FFFFFFF1FFFFFFF1FFFFFFF1FFFFFFF1FFFFFFF",
INIT_18 => X"03FFFFFF03FFFFFF03FFFFFF03FFFFFF03FFFFFF03FFFFFF03FFFFFF03FFFFFF",
INIT_19 => X"007FFFFF007FFFFF007FFFFF007FFFFF007FFFFF007FFFFF007FFFFF007FFFFF",
INIT_1a => X"000FFFFF000FFFFF000FFFFF000FFFFF000FFFFF000FFFFF000FFFFF000FFFFF",
INIT_1b => X"0001FFFF0001FFFF0001FFFF0001FFFF0001FFFF0001FFFF0001FFFF0001FFFF",
INIT_1c => X"00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF00003FFF",
INIT_1d => X"000007FF000007FF000007FF000007FF000007FF000007FF000007FF000007FF",
INIT_1e => X"000000FF000000FF000000FF000000FF000000FF000000FF000000FF000000FF",
INIT_1f => X"0000001F0000001F0000001F0000001F0000001F0000001F0000001F0000001F",
INIT_20 => X"0000000300000003000000030000000300000003000000030000000300000003",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"FFFFFFFF800000018000000180000001800000018000000180000001FFFFFFFF",
INIT_23 => X"FFFFFFFF800000018000000180000001800000018000000180000001FFFFFFFF",
INIT_24 => X"FFFFFFFF800000018000000180000001800000018000000180000001FFFFFFFF",
INIT_25 => X"FFFFFFFF800000018000000180000001800000018000000180000001FFFFFFFF",
INIT_26 => X"FFFFFFFF800000018000000180000001800000018000000180000001FFFFFFFF",
INIT_27 => X"FFFFFFFF800000018000000180000001800000018000000180000001FFFFFFFF",
INIT_28 => X"0300000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"1B60000003000000000000000000000000000000000000000000000000000000",
INIT_2a => X"1B6000001B600000030000000000000000000000000000000000000000000000",
INIT_2b => X"1B6000001B6000001B6000000300000000000000000000000000000000000000",
INIT_2c => X"1FE000001B6000001B6000001B60000003000000000000000000000000000000",
INIT_2d => X"1FEC00001FE000001B6000001B6000001B600000030000000000000000000000",
INIT_2e => X"1FFC00001FEC00001FE000001B6000001B6000001B6000000300000000000000",
INIT_2f => X"1FFC00001FEC00001FE000001B6000001B600000030000000000000000000000",
INIT_30 => X"1FFC00001FEC00001FE000001B60000003000000000000000000000000000000",
INIT_31 => X"1FEC00001FE000001B6000000300000000000000000000000000000000000000",
INIT_32 => X"1FE000001B600000030000000000000000000000000000000000000000000000",
INIT_33 => X"1B60000003000000000000000000000000000000000000000000000000000000",
INIT_34 => X"1B60000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"1B60000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"1B6000C000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"1B6006D8000000C0000000000000000000000000000000000000000000000000",
INIT_38 => X"1B6006D8000006D8000000C00000000000000000000000000000000000000000",
INIT_39 => X"1B6006D8000006D8000006D8000000C000000000000000000000000000000000",
INIT_3a => X"1B6007F8000006D8000006D8000006D8000000C0000000000000000000000000",
INIT_3b => X"1B6037F8000007F8000006D8000006D8000006D8000000C00000000000000000",
INIT_3c => X"1B603FF8000037F8000007F8000006D8000006D8000006D8000000C000000000",
INIT_3d => X"1B603FF8000037F8000007F8000006D8000006D8000000C00000000000000000",
INIT_3e => X"1B603FF8000037F8000007F8000006D8000000C0000000000000000000000000",
INIT_3f => X"1B6037F8000007F8000006D8000000C000000000000000000000000000000000")
   port map (
      DO => pixel1,      -- 1-bit Data Output
      ADDR => addres1,  -- 14-bit Address Input
      CLK => mclk,    -- Clock
      DI => "0",      -- 1-bit Data Input
      EN => '1',      -- RAM Enable Input
      SSR => '0',    -- Synchronous Set/Reset Input
      WE => '0'       -- Write Enable Input
   );  

    RAMB16_S1_inst2 : RAMB16_S1
   generic map (
      INIT => "0", --  Value of output RAM registers at startup
      SRVAL => "0", --  Ouput value upon SSR assertion
      WRITE_MODE => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
INIT_00 => X"1B6007F8000006D8000000C00000000000000000000000000000000000000000",
INIT_01 => X"1B6006D8000000C0000000000000000000000000000000000000000000000000",
INIT_02 => X"1B6006D800000000000000000000000000000000000000000000000000000000",
INIT_03 => X"1B6006D800000000000000000000000000000000000000000000000000000000",
INIT_04 => X"1B63C6D800000000000000000000000000000000000000000000000000000000",
INIT_05 => X"1B67E6D80003C000000000000000000000000000000000000000000000000000",
INIT_06 => X"1B6FF6D80007E0000003C0000000000000000000000000000000000000000000",
INIT_07 => X"1B7FFED8000FF0000007E0000003C00000000000000000000000000000000000",
INIT_08 => X"1B799ED8001FF800000FF0000007E0000003C000000000000000000000000000",
INIT_09 => X"1B799ED800199800001FF800000FF0000007E0000003C0000000000000000000",
INIT_0a => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_0b => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_0c => X"1B7FFED800199800001FF800001FF800000FF0000007E0000003C00000000000",
INIT_0d => X"1B7FFED8001FF800001FF800001FF800000FF0000007E0000003C00000000000",
INIT_0e => X"1B7FFED800199800001FF800001FF800000FF0000007E0000003C00000000000",
INIT_0f => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_10 => X"1B7FFED800199800001FF800001FF800000FF0000007E0000003C00000000000",
INIT_11 => X"1B7FFED8001FF800001FF800001FF800000FF0000007E0000003C00000000000",
INIT_12 => X"1B7FFED800199800001FF800001FF800000FF0000007E0000003C00000000000",
INIT_13 => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_14 => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_15 => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_16 => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_17 => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_18 => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_19 => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_1a => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_1b => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_1c => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_1d => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_1e => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_1f => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_20 => X"1B7FFED8001998000019F800001FF800000FF0000007E0000003C00000000000",
INIT_21 => X"1B7FFED80019F8000019F800001FF800000FF0000007E0000003C00000000000",
INIT_22 => X"1B7FFED8001998000019F800001FF800000FF0000007E0000003C00000000000",
INIT_23 => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_24 => X"1B7FFED8001998000019F800001FF800000FF0000007E0000003C00000000000",
INIT_25 => X"1B7FFED80019F8000019F800001FF800000FF0000007E0000003C00000000000",
INIT_26 => X"1B7FFED80019F8000019F800001FF800000FF0000007E0000003C00000000000",
INIT_27 => X"1B7FFED80019F8000019F800001FF800000FF0000007E0000003C00000000000",
INIT_28 => X"1B7FFED80019F8000019F800001FF800000FF0000007E0000003C00000000000",
INIT_29 => X"1B7FFED8001998000019F800001FF800000FF0000007E0000003C00000000000",
INIT_2a => X"1B7FFED800199800001FF800001FF800000FF0000007E0000003C00000000000",
INIT_2b => X"1B7FFED800199800001FF800001FF800000FF0000007E0000003C00000000000",
INIT_2c => X"1B7FFED800199800001FF800001FF800000FF0000007E0000003C00000000000",
INIT_2d => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_2e => X"1B7FFED80019980000199800001FF800000FF0000007E0000003C00000000000",
INIT_2f => X"1B7FF6D80033300000333000003FF000001FE000000FC0000007800000000000",
INIT_30 => X"1B7FE6D80066600000666000007FE000003FC000001F8000000F000000000000",
INIT_31 => X"1BFFC6D800CCC00000CCC00000FFC000007F8000003F0000001E000000000000",
INIT_32 => X"1BFF86D8019980000199800001FF800000FF0000007E0000003C000000000000",
INIT_33 => X"1BFF06D8033300000333000003FF000001FE000000FC00000078000000000000",
INIT_34 => X"1FFE06D8066600000666000007FE000003FC000001F8000000F0000000000000",
INIT_35 => X"1FFE06D8066600000666000007FE000003FC000001F8000000F0000000000000",
INIT_36 => X"1FFE06D8066600C00666000007FE000003FC000001F8000000F0000000000000",
INIT_37 => X"1FFE06D8066606D8066600C007FE000003FC000001F8000000F0000000000000",
INIT_38 => X"1FFE06D8066606D8066606D807FE00C003FC000001F8000000F0000000000000",
INIT_39 => X"1FFE37F8066606D8066606D807FE06D803FC00C001F8000000F0000000000000",
INIT_3a => X"1FFE1FF8066637F8066606D807FE06D803FC06D801F800C000F0000000000000",
INIT_3b => X"1FFE0FF006661FF8066637F807FE06D803FC06D801F806D800F000C000000000",
INIT_3c => X"1FFE1FE006663FF006666FF007FE0DB003FC0DB001F80DB000F0018000000000",
INIT_3d => X"1FFE3FC006667FE00666DFE007FE1B6003FC1B6001F81B6000F0030000000000",
INIT_3e => X"1FFE7F800666FFC00667BFC007FE36C003FC36C001F836C000F0060000000000",
INIT_3f => X"1FFE3FC006667FE00666DFE007FE1B6003FC1B6001F81B6000F0030000000000")
   port map (
      DO => pixel2,      -- 1-bit Data Output
      ADDR => addres2,  -- 14-bit Address Input
      CLK => mclk,    -- Clock
      DI => "0",      -- 1-bit Data Input
      EN => '1',      -- RAM Enable Input
      SSR => '0',    -- Synchronous Set/Reset Input
      WE => '0'       -- Write Enable Input
   );
   

   RAMB16_S1_inst3 : RAMB16_S1
   generic map (
      INIT => "0", --  Value of output RAM registers at startup
      SRVAL => "0", --  Ouput value upon SSR assertion
      WRITE_MODE => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
INIT_00 => X"1FFE1FE006663FF006666FF007FE0DB003FC0DB001F80DB000F0018000000000",
INIT_01 => X"1FFE0FF006661FF8066637F807FE06D803FC06D801F806D800F000C000000000",
INIT_02 => X"1FFE07F806660FFC06661BFC07FE036C03FC036C01F8036C00F0006000000000",
INIT_03 => X"1FFE03FC066607FE06660DFE07FE01B603FC01B601F801B600F0003000000000",
INIT_04 => X"1FFE01FE066603FF066606FF07FE00DB03FC00DB01F800DB00F0001800000000",
INIT_05 => X"1FFE03FC066607FE06660DFE07FE01B603FC01B601F801B600F0003000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"1FFE07F806660FFC06661BFC07FE036C03FC036C01F8036C00F0006000000000",
INIT_08 => X"1FFE0FF006661FF8066637F807FE06D803FC06D801F806D800F000C000000000",
INIT_09 => X"1FFE1FE006663FF006666FF007FE0DB003FC0DB001F80DB000F0018000000000",
INIT_0a => X"1FFE1FE006663FF006666FF007FE0DB003FC0DB001F80DB000F0018000000000",
INIT_0b => X"1FFE1FE006663FF006666FF007FE0DB003FC0DB001F80DB000F0018000000000",
INIT_0c => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0d => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0e => X"0000000000000000000000008000000080000000000000000000000000000000",
INIT_0f => X"00000000000000000000000080000000C0000000400000000000000000000000",
INIT_10 => X"00000000000000000000000080000000C0000000600000002000000000000000",
INIT_11 => X"00000000000000000000000080000000C0000000600000003000000010000000",
INIT_12 => X"00000000000000000000000080000000C0000000600000003800000018000000",
INIT_13 => X"00000000000000000000000080000000C0000000640000003C00000018000000",
INIT_14 => X"00000000000000000000000080000000C2000000660000003C00000018000000",
INIT_15 => X"00000000000000000000000081000000C3000000660000003C00000018000000",
INIT_16 => X"00000000000000000080000081800000C3000000660000003C00000018000000",
INIT_17 => X"000000000040000000C0000081800000C3000000660000003C00000018000000",
INIT_18 => X"002000000060000000C0000081800000C3000000660000003C00000018000000",
INIT_19 => X"003000000070000000C0000081800000C3000000660000003C00000018000000",
INIT_1a => X"003000000078000000C8000081800000C3000000660000003C00000018000000",
INIT_1b => X"003000000078000000CC000081840000C3000000660000003C00000018000000",
INIT_1c => X"003000000078000000CC000081860000C3020000660000003C00000018000000",
INIT_1d => X"003000000078000000CC000081860000C3030000660100003C00000018000000",
INIT_1e => X"003000000078000000CC000081860000C3030000660180003C00800018000000",
INIT_1f => X"003000000078000000CC000081860000C3030000660180003C00C00018004000",
INIT_20 => X"003000000078000000CC000081860000C3030000660180003C00E00018006000",
INIT_21 => X"003000000078000000CC000081860000C3030000660190003C00F00018006000",
INIT_22 => X"003000000078000000CC000081860000C3030800660198003C00F00018006000",
INIT_23 => X"003000000078000000CC000081860400C3030C00660198003C00F00018006000",
INIT_24 => X"003000000078000000CC020081860600C3030C00660198003C00F00018006000",
INIT_25 => X"003000000078010000CC030081860600C3030C00660198003C00F00018006000",
INIT_26 => X"003000800078018000CC030081860600C3030C00660198003C00F00018006000",
INIT_27 => X"003000C0007801C000CC030081860600C3030C00660198003C00F00018006000",
INIT_28 => X"003000C0007801E000CC032081860600C3030C00660198003C00F00018006000",
INIT_29 => X"003000C0007801E000CC033081860610C3030C00660198003C00F00018006000",
INIT_2a => X"003000C0007801E000CC033081860618C3030C08660198003C00F00018006000",
INIT_2b => X"003000C0007801E000CC033081860618C3030C0C660198043C00F00018006000",
INIT_2c => X"003000C0007801E000CC033081860618C3030C0C660198063C00F00218006000",
INIT_2d => X"003000C0007801E000CC033081860618C3030C0C660198063C00F00318006001",
INIT_2e => X"00180060003C00F080660198C0C3030C618186063300CC031E0078010C003000",
INIT_2f => X"000C0030801E0078C03300CC6061818630C0C303198066010F003C0006001800",
INIT_30 => X"80060018C00F003C601980663030C0C3186061810CC0330007801E0003000C00",
INIT_31 => X"C003000CE007801E300CC033181860610C3030C00660198003C00F0001800600",
INIT_32 => X"60018006F003C00F980660190C0C30300618186003300CC001E0078000C00300",
INIT_33 => X"3000C0037801E007CC03300C86061818030C0C300198066000F003C000600180",
INIT_34 => X"180060013C00F00366019806C3030C0C8186061800CC0330007801E0003000C0",
INIT_35 => X"0C0030001E0078013300CC0361818606C0C3030C80660198003C00F000180060",
INIT_36 => X"060018000F003C001980660130C0C30360618186C03300CC801E0078000C0030",
INIT_37 => X"03000C0007801E000CC03300186061813030C0C360198066C00F003C80060018",
INIT_38 => X"0180060003C00F00066019800C3030C018186061300CC033E007801EC003000C",
INIT_39 => X"00C0030001E0078003300CC0061818600C0C303098066019F003C00F60018006",
INIT_3a => X"0060018000F003C001980660030C0C3086061818CC03300C7801E0073000C003",
INIT_3b => X"003000C0007801E000CC033081860618C3030C0C660198063C00F00318006001",
INIT_3c => X"00180060003C00F080660198C0C3030C618186063300CC031E0078010C003000",
INIT_3d => X"000C0030801E0078C03300CC6061818630C0C303198066010F003C0006001800",
INIT_3e => X"80060018C00F003C601980663030C0C3186061810CC0330007801E0003000C00",
INIT_3f => X"0000000000000001000000010000000100000001000000010000000100000000")
   port map (
      DO => pixel3,      -- 1-bit Data Output
      ADDR => addres3,  -- 14-bit Address Input
      CLK => mclk,    -- Clock
      DI => "0",      -- 1-bit Data Input
      EN => '1',      -- RAM Enable Input
      SSR => '0',    -- Synchronous Set/Reset Input
      WE => '0'       -- Write Enable Input
   );
   

   RAMB16_S1_inst4 : RAMB16_S1
   generic map (
      INIT => "0", --  Value of output RAM registers at startup
      SRVAL => "0", --  Ouput value upon SSR assertion
      WRITE_MODE => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
INIT_00 => X"0000000000000003000000020000000200000002000000020000000200000000",
INIT_01 => X"0000000000000007000000040000000400000004000000040000000400000000",
INIT_02 => X"000000000000000F000000080000000800000008000000080000000800000000",
INIT_03 => X"000000000000001E000000100000001000000010000000100000001000000000",
INIT_04 => X"000000000000003D000000210000002100000021000000210000002000000000",
INIT_05 => X"000000000000007A000000420000004300000042000000420000004100000000",
INIT_06 => X"00000000000000F4000000840000008700000084000000840000008300000000",
INIT_07 => X"00000000000001E9000001090000010F00000109000001090000010600000000",
INIT_08 => X"00000000000003D2000002120000021E00000212000002120000020C00000000",
INIT_09 => X"00000000000007A5000004240000043C00000425000004250000041800000000",
INIT_0a => X"0000000000000F4B00000848000008790000084A0000084A0000083100000000",
INIT_0b => X"0000000000001E9700001090000010F300001094000010940000106300000000",
INIT_0c => X"0000000000003D2E00002121000021E60000212800002128000020C600000000",
INIT_0d => X"0000000000007A5C00004242000043CC00004250000042500000418C00000000",
INIT_0e => X"000000000000F4B90000848500008799000084A1000084A10000831900000000",
INIT_0f => X"000000000001E9730001090A00010F3200010943000109420001063300000000",
INIT_10 => X"000000000003D2E70002121400021E64000212870002128400020C6700000000",
INIT_11 => X"000000000007A5CF0004242800043CC80004250F00042508000418CF00000000",
INIT_12 => X"00000000000F4B9E000848500008799000084A1E00084A100008319E00000000",
INIT_13 => X"00000000001E973D001090A10010F3210010943D001094210010633D00000000",
INIT_14 => X"00000000003D2E7A002121420021E6420021287B002128420020C67B00000000",
INIT_15 => X"00000000007A5CF4004242840043CC85004250F70042508400418CF700000000",
INIT_16 => X"0000000000F4B9E8008485090087990A0084A1EE0084A109008319EE00000000",
INIT_17 => X"0000000001E973D101090A12010F3214010943DC01094212010633DC00000000",
INIT_18 => X"0000000003D2E7A202121424021E6428021287B802128424020C67B800000000",
INIT_19 => X"0000000007A5CF4404242848043CC85004250F70042508480418CF7000000000",
INIT_1a => X"000000000F4B9E8808485090087990A0084A1EE0084A109008319EE000000000",
INIT_1b => X"000000001E973D111090A12010F3214010943DC11094212110633DC000000000",
INIT_1c => X"000000003D2E7A232121424021E6428121287B822128424220C67B8100000000",
INIT_1d => X"000000007A5CF4474242848043CC85034250F70442508484418CF70300000000",
INIT_1e => X"00000000F4B9E88E8485090187990A0684A1EE0884A109088319EE0600000000",
INIT_1f => X"00000000E973D11C090A12020F32140C0943DC10094212100633DC0C00000000",
INIT_20 => X"00000000D2E7A239121424051E6428191287B821128424210C67B81900000000",
INIT_21 => X"00000000A5CF44722428480A3CC85032250F70432508484218CF703200000000",
INIT_22 => X"000000004B9E88E4485090147990A0644A1EE0874A109084319EE06400000000",
INIT_23 => X"00000000973D11C990A12029F32140C9943DC10F94212109633DC0C900000000",
INIT_24 => X"000000002E7A239221424052E6428192287B821E28424212C67B819200000000",
INIT_25 => X"000000005CF44724428480A5CC85032550F7043D508484258CF7032400000000",
INIT_26 => X"00000000B9E88E498509014A990A064AA1EE087AA109084A19EE064900000000",
INIT_27 => X"0000000073D11C930A12029432140C9443DC10F44212109433DC0C9300000000",
INIT_28 => X"00000000E7A23926142405296428192987B821E98424212967B8192600000000",
INIT_29 => X"00000000CF44724C28480A52C85032520F7043D208484252CF70324C00000000",
INIT_2a => X"000000009E88E498509014A490A064A51EE087A5109084A59EE0649900000000",
INIT_2b => X"000000003D11C930A12029492140C94A3DC10F4A2121094A3DC0C93200000000",
INIT_2c => X"000000007A23926142405292428192947B821E94424212947B81926400000000",
INIT_2d => X"00000000F44724C28480A52585032529F7043D2984842529F70324C900000000",
INIT_2e => X"00000000E88E498509014A4A0A064A52EE087A5209084A52EE06499200000000",
INIT_2f => X"00000000D11C930A12029495140C94A4DC10F4A4121094A4DC0C932400000000",
INIT_30 => X"00000000A23926142405292A28192949B821E94924212949B819264900000000",
INIT_31 => X"0000000044724C28480A5254503252927043D2924842529270324C9200000000",
INIT_32 => X"0000000088E498509014A4A8A064A524E087A5249084A524E064992400000000",
INIT_33 => X"0000000011C930A02029495040C94A48C10F4A4821094A48C0C9324800000000",
INIT_34 => X"0000000023926140405292A081929490821E9490421294908192649000000000",
INIT_35 => X"000000004724C28080A5254003252920043D2920842529200324C92000000000",
INIT_36 => X"000000008E498500014A4A80064A5240087A5240084A52400649924000000000",
INIT_37 => X"000000001C930A00029495000C94A48010F4A4801094A4800C93248000000000",
INIT_38 => X"000000003926140005292A001929490021E94900212949001926490000000000",
INIT_39 => X"00000000724C28000A5254003252920043D2920042529200324C920000000000",
INIT_3a => X"00000000E498500014A4A80064A5240087A5240084A524006499240000000000",
INIT_3b => X"00000000C930A00029495000C94A48000F4A4800094A4800C932480000000000",
INIT_3c => X"00000000926140005292A000929490001E949000129490009264900000000000",
INIT_3d => X"0000000024C28000A5254000252920003D2920002529200024C9200000000000",
INIT_3e => X"00000000498500004A4A80004A5240007A5240004A5240004992400000000000",
INIT_3f => X"00000000930A00009495000094A48000F4A4800094A480009324800000000000")
   port map (
      DO => pixel4,      -- 1-bit Data Output
      ADDR => addres4,  -- 14-bit Address Input
      CLK => mclk,    -- Clock
      DI => "0",      -- 1-bit Data Input
      EN => '1',      -- RAM Enable Input
      SSR => '0',    -- Synchronous Set/Reset Input
      WE => '0'       -- Write Enable Input
   );
   


end Behavioral;
