------------------------------------------------------------------------
--	OscillatorsUnit.vhd
------------------------------------------------------------------------
--	Author:	Lucian Chetan
------------------------------------------------------------------------
--	Software version: Xilinx WebPack ISE 8.1i
------------------------------------------------------------------------
--	This module groups the modules that:
--		-	generates the notes periods that the oscillators will use ("NoteMemory"),
--		-	generates the four waves according to the four note periods ("OscillatorGroup"),
--		-	resample the data at a constant 48 kHz ("Sampler").
------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity OscillatorsUnit is
	port (
		clk					: in STD_LOGIC; -- Master clock (50 MHz)
		rst					: in STD_LOGIC; -- Reset button (synchronous reset)
		waveType				: in STD_LOGIC; -- The type of wave generated by the oscillators: '0' = sawtooth, '1'  = square
		oscillatorStatus	: in STD_LOGIC_VECTOR(3 downto 0); -- The status of the 4 oscillators
		noteAddress0		: in STD_LOGIC_VECTOR(4 downto 0); -- The note handled by the first oscillator
		noteAddress1		: in STD_LOGIC_VECTOR(4 downto 0); -- The note handled by the second oscillator
		noteAddress2		: in STD_LOGIC_VECTOR(4 downto 0); -- The note handled by the third oscillator
		noteAddress3		: in STD_LOGIC_VECTOR(4 downto 0); -- The note handled by the fourth oscillator
		outputWave			: out STD_LOGIC_VECTOR(7 downto 0) -- The resulting wave
	);
end OscillatorsUnit;

architecture Behavioral of OscillatorsUnit is

	-- This component represents the memory of note periods.
	component NoteMemory is
		port (
			noteAddress0	: in STD_LOGIC_VECTOR(4 downto 0);
			noteAddress1	: in STD_LOGIC_VECTOR(4 downto 0);
			noteAddress2	: in STD_LOGIC_VECTOR(4 downto 0);
			noteAddress3	: in STD_LOGIC_VECTOR(4 downto 0);
			notePeriod0		: out STD_LOGIC_VECTOR(10 downto 0);
			notePeriod1		: out STD_LOGIC_VECTOR(10 downto 0);
			notePeriod2		: out STD_LOGIC_VECTOR(10 downto 0);
			notePeriod3		: out STD_LOGIC_VECTOR(10 downto 0)
		);
	end component;

	-- This component represents the 4 oscillators which, if enabled, oscillate according to the note period.
	component OscillatorGroup is
		port (
			clk					: in STD_LOGIC;
			rst					: in STD_LOGIC;
			waveType				: in STD_LOGIC;
			oscillatorStatus	: in STD_LOGIC_VECTOR(3 downto 0);
			notePeriod0			: in STD_LOGIC_VECTOR(10 downto 0);
			notePeriod1			: in STD_LOGIC_VECTOR(10 downto 0);
			notePeriod2			: in STD_LOGIC_VECTOR(10 downto 0);
			notePeriod3			: in STD_LOGIC_VECTOR(10 downto 0);
			outputWave			: out STD_LOGIC_VECTOR(7 downto 0)
		);
	end component;

	-- This component samples at 48 kHz the data generated by the oscillators.
	component Sampler is
		port (
			clk		: in STD_LOGIC;
			dataIn	: in STD_LOGIC_VECTOR(7 downto 0);
			dataOut	: out STD_LOGIC_VECTOR(7 downto 0)
		);
	end component;

	signal notePeriod0		: STD_LOGIC_VECTOR(10 downto 0);
	signal notePeriod1		: STD_LOGIC_VECTOR(10 downto 0);
	signal notePeriod2		: STD_LOGIC_VECTOR(10 downto 0);
	signal notePeriod3		: STD_LOGIC_VECTOR(10 downto 0);
	signal outputWave_temp	: STD_LOGIC_VECTOR(7 downto 0);

begin

	NoteMemory_Map: NoteMemory port map (
		noteAddress0 => noteAddress0,
		noteAddress1 => noteAddress1,
		noteAddress2 => noteAddress2,
		noteAddress3 => noteAddress3,
		notePeriod0 => notePeriod0,
		notePeriod1 => notePeriod1,
		notePeriod2 => notePeriod2,
		notePeriod3 => notePeriod3
	);

	OscillatorGroup_Map: OscillatorGroup port map (
		clk => clk,
		rst => rst,
		waveType => waveType,
		oscillatorStatus => oscillatorStatus,
		notePeriod0 => notePeriod0,
		notePeriod1 => notePeriod1,
		notePeriod2 => notePeriod2,
		notePeriod3 => notePeriod3,
		outputWave => outputWave_temp
	);

	Sampler_Map: Sampler port map (
		clk => clk,
		dataIn => outputWave_temp,
		dataOut => outputWave
	);

end Behavioral;