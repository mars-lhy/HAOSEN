
-------------------------------------------------------------------------------
--     ChMap.vhd -- Stores 8x8 pixel patterns for the basic characters
-------------------------------------------------------------------------------
--		Inputs:
--			Ascii(5:0)	The predefined code of the actual character
--			Line(2:0)	Number of the  pixel line from the previously defined char
--		Outputs:
--			Data(7:0)	The pixel codes of the character line: ROM(Ascii&Line)
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--  Uncomment the following lines to use the declarations that are
--  provided for instantiating Xilinx primitive components.
--library UNISIM;
--use UNISIM.VComponents.all;

entity chmap is
    Port ( ascii : in std_logic_vector(5 downto 0);
           line : in std_logic_vector(2 downto 0);
           data : out std_logic_vector(7 downto 0));
end chmap;

architecture Behavioral of chmap is
	type ROM_Array is array (0 to 511)
		of std_logic_vector(7 downto 0);

	constant Content: ROM_Array := (
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00111000",--A
		"01000100",
		"01000100",
		"01000100",
		"01111100",
		"01000100",
		"01000100",
		"00000000",
		"01111000",--B
		"01000100",
		"01000100",
		"01111000",
		"01000100",
		"01000100",
		"01111000",
		"00000000",
		"00111000",--C
		"01000100",
		"01000000",
		"01000000",
		"01000000",
		"01000100",
		"00111000",
		"00000000",
		"01110000",--D
		"01001000",
		"01000100",
		"01000100",
		"01000100",
		"01001000",
		"01110000",
		"00000000",
		"01111100",--E
		"01000000",
		"01000000",
		"01111000",
		"01000000",
		"01000000",
		"01111100",
		"00000000",
		"01111100",--F
		"01000000",
		"01000000",
		"01111000",
		"01000000",
		"01000000",
		"01000000",
		"00000000",
		"00111000",--G
		"01000100",
		"01000000",
		"01011100",
		"01000100",
		"01000100",
		"00111000",
		"00000000",
		"01000100",--H
		"01000100",
		"01000100",
		"01111100",
		"01000100",
		"01000100",
		"01000100",
		"00000000",
		"00111000",--I
		"00010000",
		"00010000",
		"00010000",
		"00010000",
		"00010000",
		"00111000",
		"00000000",
		"00011100",--J
		"00001000",
		"00001000",
		"00001000",
		"00001000",
		"00101000",
		"00110000",
		"00000000",
		"01000100",--K
		"01001000",
		"01010000",
		"01100000",
		"01010000",
		"01001000",
		"01000100",
		"00000000",
		"01000000",--L
		"01000000",
		"01000000",
		"01000000",
		"01000000",
		"01000000",
		"01111100",
		"00000000",
		"01000100",--M
		"01101100",
		"01010100",
		"01000100",
		"01000100",
		"01000100",
		"00000000",
		"00000000",
		"01000100",--N
		"01000100",
		"01100100",
		"01010100",
		"01001100",
		"01000100",
		"00000000",
		"00000000",
		"00111000",--O
		"01000100",
		"01000100",
		"01000100",
		"01000100",
		"01000100",
		"00111000",
		"00000000",
		"01111000",--P
		"01000100",
		"01000100",
		"01111000",
		"01000000",
		"01000000",
		"01000000",
		"00000000",
		"00111000",--Q
		"01000100",
		"01000100",
		"01000100",
		"01010100",
		"01001000",
		"00110100",
		"00000000",
		"01111000",--R
		"01000100",
		"01000100",
		"01111000",
		"01010000",
		"01001000",
		"01000100",
		"00000000",
		"00111100",--S
		"01000000",
		"01000000",
		"00111000",
		"00000100",
		"00000100",
		"01111000",
		"00000000",
		"01111100",--T
		"00010000",
		"00010000",
		"00010000",
		"00010000",
		"00010000",
		"00010000",
		"00000000",
		"01000100",--U
		"01000100",
		"01000100",
		"01000100",
		"01000100",
		"01000100",
		"00111000",
		"00000000",
		"01000100",--V
		"01000100",
		"01000100",
		"01000100",
		"01000100",
		"00101000",
		"00010000",
		"00000000",
		"01000100",--W
		"01000100",
		"01000100",
		"01010100",
		"01010100",
		"01010100",
		"00101000",
		"00000000",
		"01000100",--X
		"01000100",
		"00101000",
		"00010000",
		"00101000",
		"01000100",
		"01000100",
		"00000000",
		"01000100",--Y
		"01000100",
		"01000100",
		"00101000",
		"00010000",
		"00010000",
		"00010000",
		"00000000",
		"01111100",--Z
		"00000100",
		"00001000",
		"00010000",
		"00100000",
		"01000000",
		"01111100",
		"00000000",
		"00111000",--O
		"01000100",
		"01001100",
		"01010100",
		"01100100",
		"01000100",
		"00111000",
		"00000000",
		"00010000",--1
		"00110000",
		"00010000",
		"00010000",
		"00010000",
		"00010000",
		"00111000",
		"00000000",
		"00111000",--2
		"01000100",
		"00000100",
		"00001000",
		"00010000",
		"00100000",
		"01111100",
		"00000000",
		"01111100",--3
		"01001000",
		"00010000",
		"00001000",
		"00000100",
		"01000100",
		"00111000",
		"00000000",
		"00001000",--4
		"00011000",
		"00101000",
		"01001000",
		"01111100",
		"00001000",
		"00001000",
		"00000000",
		"01111100",--5
		"01000000",
		"01111000",
		"00000100",
		"00000100",
		"01000100",
		"00111000",
		"00000000",
		"00011000",--6
		"00100000",
		"01000000",
		"01111000",
		"01000100",
		"01000100",
		"00111000",
		"00000000",
		"01111100",--7
		"00000100",
		"00001000",
		"00010000",
		"00100000",
		"00100000",
		"00100000",
		"00000000",
		"00111000",--8
		"01000100",
		"01000100",
		"00111000",
		"01000100",
		"01000100",
		"00111000",
		"00000000",
		"00111000",--9
		"01000100",
		"01000100",
		"00111000",
		"00000100",
		"00000100",
		"00110000",
		"00000000",
		"00000000",--space
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",--,
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00110000",
		"00010000",
		"00100000",
		"00000000",--.
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00110000",
		"00110000",
		"00000000",
		"00000000",--/
		"00000100",
		"00001000",
		"00010000",
		"00100000",
		"01000000",
		"00000000",
		"00000000",
		"00000000",--;
		"00110000",
		"00110000",
		"00000000",
		"00000000",
		"00110000",
		"00010000",
		"00100000",
		"00110000",--'
		"00010000",
		"00100000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",--\
		"01000000",
		"00100000",
		"00010000",
		"00001000",
		"00000100",
		"00000000",
		"00000000",
		"00111000",--[
		"00100000",
		"00100000",
		"00100000",
		"00100000",
		"00100000",
		"00111000",
		"00000000",
		"00111000",--]
		"00001000",
		"00001000",
		"00001000",
		"00001000",
		"00001000",
		"00111000",
		"00000000",
		"00000000",---
		"00000000",
		"00000000",
		"01111100",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",--=
		"00000000",
		"01111100",
		"00000000",
		"01111100",
		"00000000",
		"00000000",
		"00000000",
		"00100000",--`
		"00010000",
		"00001000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		OTHERS => "00000000");

	signal addr : std_logic_vector(8 downto 0) := "000000000";

begin
	
	addr(8 downto 0) <= ascii(5 downto 0) & line(2 downto 0);
	data <= Content(conv_integer(addr)); 
	
end Behavioral;
