------------------------------------------------------------------------
--	CircularMemory.vhd
------------------------------------------------------------------------
--	Author:	Digilent
--				Lucian Chetan (modified state machine)
------------------------------------------------------------------------
--	Software version:	Xilinx WebPack ISE 8.1i
------------------------------------------------------------------------
--	This module represents a 16384 x 8-bit memory that stores the samples
--	generated by the oscillators. The time difference between two consecutive
--	addresses is 1 / 48 kHz ~= 20 us. The time difference between the oldest
--	sample and the newest sample is 16383 * 20 us = 16383 / 48 kHz = 0,341 seconds.
------------------------------------------------------------------------

library ieee;
use ieee.STD_LOGIC_1164.all;
use ieee.STD_LOGIC_unsigned.all;

entity CircularMemory is
	port (
		clk		: in STD_LOGIC; -- Master clock (50 MHz)
		we			: in STD_LOGIC; -- Write enable
		address	: in STD_LOGIC_VECTOR(13 downto 0); -- Write/read address
		dataIn	: in STD_LOGIC_VECTOR(7 downto 0); -- Write data
		dataOut	: out STD_LOGIC_VECTOR(7 downto 0) -- Read data
	);
end CircularMemory;

architecture Behavioral of CircularMemory is

	signal readAddress: STD_LOGIC_VECTOR(13 downto 0);

	-- Memory size is 16384 bytes, in order to accomodate delays large enough for the 'delay' and 'echo' effects.
	-- Maximum delay is 16383 * 20 us = 327,66 ms.
	type ram_type is array (0 to 16383) of STD_LOGIC_VECTOR (7 downto 0);
	signal RAM: ram_type;

begin
	process (clk)
	begin
		if rising_edge(clk) then
			if (we = '1') then
				RAM(conv_integer(address)) <= dataIn;
			end if;
			readAddress <= address;
		end if;
	end process;
	
	dataOut <= RAM(conv_integer(readAddress));
	
end Behavioral;