------------------------------------------------------------------------
--	UsbUnit.vhd
------------------------------------------------------------------------
--	Author:	Digilent
--				Lucian Chetan (modified state machine)
------------------------------------------------------------------------
--	Software version:	Xilinx WebPack ISE 8.1i
------------------------------------------------------------------------
--	This module implements the state machine described in the Digilent
--	Parallel Interface Model, with few modifications.
--	There are one address register and nine data registers. Their purpose is
--	to store the notes that the PC sends for playing on the FPGA board,
--	control the effects and the voice that the oscillators generate.
------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity UsbUnit is
	port (
		clk				: in STD_LOGIC; -- Master clock (50 MHz)
		eppAstb			: in STD_LOGIC; -- EPP protocol address strobe
		eppDstb			: in STD_LOGIC; -- EPP protocol data strobe
		eppWrite			: in STD_LOGIC; -- EPP protocol write strobe
		eppWait			: out STD_LOGIC; -- EPP protocol wait strobe
		eppDataBus		: inout STD_LOGIC_VECTOR(7 downto 0); -- EPP protocol data lines

		midiDirection	: in STD_LOGIC; -- Direction of MIDI messages: 0 = board -> PC/board; 1 = PC -> board
		midiNote0		: in STD_LOGIC_VECTOR(4 downto 0); -- The first note generated by the keyboard
		midiNote1		: in STD_LOGIC_VECTOR(4 downto 0); -- The second note generated by the keyboard
		midiNote2		: in STD_LOGIC_VECTOR(4 downto 0); -- The third note generated by the keyboard
		midiNote3		: in STD_LOGIC_VECTOR(4 downto 0); -- The fourth note generated by the keyboard
		midiStatus		: in STD_LOGIC_VECTOR(3 downto 0); -- The status generated by the keyboard

		usbNote0			: out STD_LOGIC_VECTOR(4 downto 0); -- The first note received from the PC
		usbNote1			: out STD_LOGIC_VECTOR(4 downto 0); -- The second note received from the PC
		usbNote2			: out STD_LOGIC_VECTOR(4 downto 0); -- The third note received from the PC
		usbNote3			: out STD_LOGIC_VECTOR(4 downto 0); -- The fourth note received from the PC
		usbStatus		: out STD_LOGIC_VECTOR(3 downto 0); -- The status received from the PC

		control			: out STD_LOGIC_VECTOR(7 downto 0); -- Register that controls the MIDI directin, oscillator voice and effect selection
		parameter0		: out STD_LOGIC_VECTOR(7 downto 0); -- Register that controls the effects
		parameter1		: out STD_LOGIC_VECTOR(7 downto 0); -- Feedback value register
		parameter2		: out STD_LOGIC_VECTOR(7 downto 0); -- Wet value register
		parameter3		: out STD_LOGIC_VECTOR(7 downto 0) -- Dry value register
	);
end UsbUnit;

architecture Behavioral of UsbUnit is

	type states is (ready, addressWrite1, addressWrite2, addressRead1,
		addressRead2, dataWrite1, dataWrite2, dataRead1, dataRead2);
	signal currentState, nextState: states;

	signal eppDir		: STD_LOGIC;
	signal eppAwr		: STD_LOGIC;
	signal eppDwr		: STD_LOGIC;
	signal eppBusOut	: STD_LOGIC_VECTOR(7 downto 0);
	signal eppBusIn	: STD_LOGIC_VECTOR(7 downto 0);
	signal regEppAddr	: STD_LOGIC_VECTOR(7 downto 0);
	signal regNote0	: STD_LOGIC_VECTOR(7 downto 0);
	signal regNote1	: STD_LOGIC_VECTOR(7 downto 0);
	signal regNote2	: STD_LOGIC_VECTOR(7 downto 0);
	signal regNote3	: STD_LOGIC_VECTOR(7 downto 0);
	signal regControl	: STD_LOGIC_VECTOR(7 downto 0);
	signal regParam0	: STD_LOGIC_VECTOR(7 downto 0);
	signal regParam1	: STD_LOGIC_VECTOR(7 downto 0); -- The "feedback" register
	signal regParam2	: STD_LOGIC_VECTOR(7 downto 0); -- The "wet" register
	signal regParam3	: STD_LOGIC_VECTOR(7 downto 0) := x"FF"; -- The "dry" register (at power-up it must be x"FF")

begin

	eppBusIn <= eppDataBus; -- the input data bus receives the data bus value
	eppDataBus <= eppBusOut when (eppWrite = '1' and eppDir = '1') else "ZZZZZZZZ"; -- the data bus value receives the value of the output bus only during read cycles
	eppBusOut <= -- the selected register outputs its value on the output bus
		regControl when (regEppAddr = x"00") else
		regNote0 when (regEppAddr = x"01") else
		regNote1 when (regEppAddr = x"02") else
		regNote2 when (regEppAddr = x"03") else
		regNote3 when (regEppAddr = x"04") else
		regParam0 when (regEppAddr = x"80") else
		regParam1 when (regEppAddr = x"81") else
		regParam2 when (regEppAddr = x"82") else
		regParam3 when (regEppAddr = x"83") else
		"00000000";

	control <= regControl;
	parameter0 <= regParam0;
	parameter1 <= regParam1;
	parameter2 <= regParam2;
	parameter3 <= regParam3;

	eppWait <=
		'1' when ((currentState = addressWrite2) or
				(currentState = addressRead2) or
				(currentState = dataWrite2) or
				(currentState = dataRead2)) else
		'0';
	eppDir <=
		'1' when ((currentState = addressRead1) or
				(currentState = addressRead2) or
				(currentState = dataRead1) or
				(currentState = dataRead2)) else
		'0';
	eppAwr <= '1' when (currentState = addressWrite1) else '0';
	eppDwr <= '1' when (currentState = dataWrite1) else '0';


	state_transition: process (clk)
	begin
		if rising_edge(clk) then
			currentState <= nextState;
		end if;
	end process;


	state_machine: process (currentState, nextState, eppAstb, eppDstb, eppWrite)
	begin
		case currentState is
			when ready =>
				if (eppAstb = '0' and eppWrite = '0') then
					nextState <= addressWrite1;
				elsif (eppAstb = '0' and eppWrite = '1') then
					nextState <= addressRead1;
				elsif (eppDstb = '0' and eppWrite = '0') then
					nextState <= dataWrite1;
				elsif (eppDstb = '0' and eppWrite = '1') then
					nextState <= dataRead1;
				else
					nextState <= ready; -- if both strobes are '1', stay in the current state
				end if;

			when addressWrite1 =>
				nextState <= addressWrite2;

			when addressWrite2 =>
				-- waiting for the host to output '1' on the address strobe
				if (eppAstb = '0') then
					nextState <= addressWrite2;
				else
					nextState <= ready;
				end if;

			when addressRead1 =>
				nextState <= addressRead2;

			when addressRead2 =>
				-- waiting for the host to output '1' on the address strobe
				if (eppAstb = '0') then
					nextState <= addressRead2;
				else
					nextState <= ready;
				end if;

			when dataWrite1 =>
				nextState <= dataWrite2;

			when dataWrite2 =>
				-- waiting for the host to output '1' on the data strobe
				if (eppDstb = '0') then
					nextState <= dataWrite2;
				else
					nextState <= ready;
				end if;

			when dataRead1 =>
				nextState <= dataRead2;

			when dataRead2 =>
				-- waiting for the host to output '1' on the data strobe
				if (eppDstb = '0') then
					nextState <= dataRead2;
				else
					nextState <= ready;
				end if;

			when others =>
				nextState <= ready;

		end case;
	end process;


	write_address_register: process (clk)
	begin
		if rising_edge(clk) then
			if (eppAwr = '1') then
				regEppAddr <= eppBusIn;
			end if;
		end if;
	end process;


	write_control_register: process (clk)
	begin
		if rising_edge(clk) then
			if (eppDwr = '1' and regEppAddr = x"00") then
				regControl <= eppBusIn;
			end if;
		end if;
	end process;


	write_param0_register: process (clk)
	begin
		if rising_edge(clk) then
			if (eppDwr = '1' and regEppAddr = x"80") then
				regParam0 <= eppBusIn;
			end if;
		end if;
	end process;


	write_param1_register: process (clk)
	begin
		if rising_edge(clk) then
			if (eppDwr = '1' and regEppAddr = x"81") then
				regParam1 <= eppBusIn;
			end if;
		end if;
	end process;


	write_param2_register: process (clk)
	begin
		if rising_edge(clk) then
			if (eppDwr = '1' and regEppAddr = x"82") then
				regParam2 <= eppBusIn;
			end if;
		end if;
	end process;


	write_param3_register: process (clk)
	begin
		if rising_edge(clk) then
			if (eppDwr = '1' and regEppAddr = x"83") then
				regParam3 <= eppBusIn;
			end if;
		end if;
	end process;


	store_notes: process (clk)
	begin
		if rising_edge(clk) then
			if (midiDirection = '1') then
				usbNote0 <= regNote0(4 downto 0);
				usbNote1 <= regNote1(4 downto 0);
				usbNote2 <= regNote2(4 downto 0);
				usbNote3 <= regNote3(4 downto 0);
				usbStatus(0) <= regNote0(7);
				usbStatus(1) <= regNote1(7);
				usbStatus(2) <= regNote2(7);
				usbStatus(3) <= regNote3(7);
			end if;
		end if;
	end process;


	write_note0_register: process (clk)
	begin
		if rising_edge(clk) then
			if (midiDirection = '1') then -- the PC sends data in order to play a MIDI file on the board
				if (eppDwr = '1' and regEppAddr = x"01") then
					regNote0 <= eppBusIn;
				end if;
			else -- the board sends data to PC in order to record a MIDI file
				regNote0 <= midiStatus(0) & "00" & midiNote0;
			end if;
		end if;
	end process;


	write_note1_register: process (clk)
	begin
		if rising_edge(clk) then
			if (midiDirection = '1') then
				if (eppDwr = '1' and regEppAddr = x"02") then
					regNote1 <= eppBusIn;
				end if;
			else
				regNote1 <= midiStatus(1) & "00" & midiNote1;
			end if;
		end if;
	end process;


	write_note2_register: process (clk)
	begin
		if rising_edge(clk) then
			if (midiDirection = '1') then
				if (eppDwr = '1' and regEppAddr = x"03") then
					regNote2 <= eppBusIn;
				end if;
			else
				regNote2 <= midiStatus(2) & "00" & midiNote2;
			end if;
		end if;
	end process;


	write_note3_register: process (clk)
	begin
		if rising_edge(clk) then
			if (midiDirection = '1') then
				if (eppDwr = '1' and regEppAddr = x"04") then
					regNote3 <= eppBusIn;
				end if;
			else
				regNote3 <= midiStatus(3) & "00" & midiNote3;
			end if;
		end if;
	end process;

end Behavioral;