------------------------------------------------------------------------
--	Oscillator.vhd
------------------------------------------------------------------------
--	Author:	Lucian Chetan
------------------------------------------------------------------------
--	Software version: Xilinx WebPack ISE 8.1i
------------------------------------------------------------------------
--	This module groups the modules that:
--		-	generate a basic wave according to the note period ("BasicOscillator"),
--		-	modulate the basic wave using the ADSR envelope model ("Enveloper").
------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Oscillator is
	port (
		clk					: in STD_LOGIC; -- Master clock (50 MHz)
		rst					: in STD_LOGIC; -- Reset button (synchronous reset)
		waveType				: in STD_LOGIC; -- The type of wave generated by the oscillator: '0' = sawtooth, '1'  = square
		oscillatorStatus	: in STD_LOGIC; -- The status of the oscillator
		notePeriod			: in STD_LOGIC_VECTOR(10 downto 0); -- The period of the note
		outputWave			: out STD_LOGIC_VECTOR(15 downto 0) -- The generated wave
	);
end Oscillator;

architecture Behavioral of Oscillator is

	-- This component represents the oscillator that generates a basic waveform, according to the period
	component BasicOscillator is
		port (
			clk				: in STD_LOGIC;
			rst				: in STD_LOGIC;
			waveType			: in STD_LOGIC;
			changePeriod	: in STD_LOGIC;
			period			: in STD_LOGIC_VECTOR(10 downto 0);
			basicWave		: out STD_LOGIC_VECTOR(7 downto 0)
		);
	end component;
	
	-- This component generates an amplitude modulated wave, using the ADSR model.
	component Enveloper is
		port (
			clk					: in STD_LOGIC;
			rst					: in STD_LOGIC;
			oscillatorStatus	: in STD_LOGIC;
			basicWave			: in STD_LOGIC_VECTOR(7 downto 0);
			envelopeIdle		: out STD_LOGIC;
			modulatedWave		: out STD_LOGIC_VECTOR(15 downto 0)
		);
	end component;
	
	signal envelopeIdle	: STD_LOGIC;
	signal basicWave_temp	: STD_LOGIC_VECTOR(7 downto 0);

begin

	BasicOscillator_Map: BasicOscillator port map (
		clk => clk,
		rst => rst,
		waveType => waveType,
		changePeriod => envelopeIdle,
		period => notePeriod,
		basicWave => basicWave_temp
	);
	
	Enveloper_Map: Enveloper port map (
		clk => clk,
		rst => rst,
		oscillatorStatus => oscillatorStatus,
		basicWave => basicWave_temp,
		envelopeIdle => envelopeIdle,
		modulatedWave => outputWave
	);

end Behavioral;