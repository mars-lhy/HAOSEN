------------------------------------------------------------------------
--	Adder.vhd
------------------------------------------------------------------------
--	Author:	Lucian Chetan
------------------------------------------------------------------------
--	Software version: Xilinx WebPack ISE 8.1i
------------------------------------------------------------------------
--	This module adds four 16-bit values and divides the result by 256.
--	The module takes as inputs the waves generated by the oscillators after
--	being modulated in amplitude (multiplied by values between 0 and 256).
--	Dividing by 256 is necessary in order to obtain the 8-bit values that
--	will be sent to the digital-to-analog converter.
------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Adder is
	port (
		a, b, c, d: in std_logic_vector(15 downto 0);
		output: out std_logic_vector(7 downto 0)
	);
end Adder;

architecture Behavioral of Adder is

	signal sum: std_logic_vector(15 downto 0);
	
begin

	sum <= a + b + c + d;
	output <= sum(15 downto 8); -- division by 256
	
end Behavioral;