------------------------------------------------------------------------
-- pixel_clock_switcher.vhd
------------------------------------------------------------------------
-- Author : Ulrich Zolt�n
--          Copyright 2006 Digilent, Inc.
------------------------------------------------------------------------
-- Software version : Xilinx ISE 7.1.04i
--                    WebPack
-- Device	        : 3s200ft256-4
------------------------------------------------------------------------
-- This file contains the logic to switch the pixel clock used,
-- depending on the resolution.
------------------------------------------------------------------------
--  Behavioral description
------------------------------------------------------------------------
-- Uses a BUFGMUX device primitive to switch between input pixel clocks,
-- generated by DCMs, the select line being the resolution input. The
-- output of this device primitive is placed on a global clock line,
-- to minimize skew.
-- Clock switching is a pretentious process, and if not done, with
-- BUFGMUX, the logic might not work as intended.
------------------------------------------------------------------------
--  Port definitions
------------------------------------------------------------------------
-- pixel_clk_25MHz   - input pin, from dcm_25MHz
--                   - the 640x480 pixel clock, that runs at 25MHz
-- pixel_clk_40MHz   - input pin, from dcm_40MHz
--                   - the 800x600 pixel clock, that runs at 40MHz
-- resolution        - input pin, from resolution_switcher
--                   - indicates with clock to choose
--                   - pixel_clk_25MHz when resolution = '0'
--                   - pixel_clk_40MHz when resolution = '1'
-- pixel_clk         - output pin
--                   - the selected pixel clock
------------------------------------------------------------------------
-- Revision History:
-- 09/18/2006(UlrichZ): created
------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- simulation library
library UNISIM;
use UNISIM.VComponents.all;

-- the pixel_clock_switcher entity declaration
-- read above for behavioral description and port definitions.
entity pixel_clock_switcher is
port(
   pixel_clk_25MHz   : in std_logic;
   pixel_clk_40MHz   : in std_logic;
   resolution        : in std_logic;
   pixel_clk         : out std_logic
);
end pixel_clock_switcher;

architecture Behavioral of pixel_clock_switcher is

begin

   -- instantiate a BUFGMUX device primitive that
   -- has inputs the 2 pixel clock generated by the
   -- DCMs and has as select line the resolution.
   -- This way pixel_clk_25MHz will be selected
   -- when resolution is '0', else pixel_clk_40MHz
   -- The output of the BUFGMUX (pixel_clk) is using
   -- a global clock line.
   BUFGMUX_inst : BUFGMUX
   port map (
      O => pixel_clk,         -- Clock MUX output
      I0 => pixel_clk_25MHz,  -- Clock0 input
      I1 => pixel_clk_40MHz,  -- Clock1 input
      S => resolution         -- Clock select input
   );

end Behavioral;