------------------------------------------------------------------------
--	BasicOscillator.vhd
------------------------------------------------------------------------
--	Author:	Lucian Chetan
------------------------------------------------------------------------
--	Software version: Xilinx WebPack ISE 8.1i
------------------------------------------------------------------------
--	This module generates the basic wave according to the note period.
--	It is capable of generating sawtooth waves which are obtained by
--	simply counting from 0 to 255, and square waves which are obtained
--	by comparing the sawtooth wave with the threshold value of 128.
------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity BasicOscillator is
	port (
		clk				: in STD_LOGIC; -- Master clock (50 MHz)
		rst				: in STD_LOGIC; -- Reset button (synchronous reset)
		waveType			: in STD_LOGIC; -- The type of wave generated by the oscillator: '0' = sawtooth, '1'  = square
		changePeriod	: in STD_LOGIC; -- Flag that determines the period to change only when the ADSR process is idle
		period			: in STD_LOGIC_VECTOR(10 downto 0); -- The period corresponding to the note
		basicWave		: out STD_LOGIC_VECTOR(7 downto 0) -- The generated wave
	);
end BasicOscillator;

architecture Behavioral of BasicOscillator is

	signal counter				: STD_LOGIC_VECTOR(16 downto 0);
	signal value				: STD_LOGIC_VECTOR(7 downto 0);
	signal period_temp		: STD_LOGIC_VECTOR(10 downto 0);
	signal sawtooth, square	: STD_LOGIC_VECTOR(7 downto 0);

begin

	-- This process reads the period only when the ADSR enveloping process is idle.
	-- This prevents period change during note playing.
	process (clk)
	begin
		if rising_edge(clk) then
			if (changePeriod = '1') then
				period_temp <= period;
			end if;
		end if;
	end process;


	-- This process counts from 0 to 255 using the note period.
	process (clk)
	begin
		if rising_edge(clk) then
			if (rst = '1') then
				counter <= (others => '0');
				value <= (others => '0');
			else
				if (counter < period_temp) then
					counter <= counter + 1;
				else
					counter <= (others => '0');
					value <= value + 1; -- The sawtooth value is increased at the end of the period. (256 increments require a period 256 times smaller so that the note has the right frequency.)
				end if;
			end if;
		end if;
	end process;


	sawtooth <= value;
	square <=
		x"00" when (value < 128) else
		x"FF";
	basicWave <= -- The 'basicWave' signal outputs the sawtooth or square wave
		sawtooth when (waveType = '0') else
		square;

end Behavioral;